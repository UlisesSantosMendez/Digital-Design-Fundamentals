module numeros ( 
	x,
	f
	) ;

input [0:3] x;
inout  f;
