module codificador ( 
	a_IBV,
	d
	) ;

input [3:0] a_IBV;
inout [3:0] d;
