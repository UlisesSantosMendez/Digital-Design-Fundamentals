module registro ( 
	r,
	er,
	clk,
	reg
	) ;

input [3:0] r;
input  er;
input  clk;
inout [3:0] reg;
