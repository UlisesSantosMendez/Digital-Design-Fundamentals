module rs ( 
	s,
	r,
	clk,
	q,
	qn
	) ;

input  s;
input  r;
input  clk;
inout  q;
inout  qn;
