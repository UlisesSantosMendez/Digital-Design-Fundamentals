module contador ( 
	sum,
	sensor,
	reset,
	compara,
	q
	) ;

inout [7:0] sum;
input  sensor;
input  reset;
inout [7:0] compara;
inout [7:0] q;
