module d ( 
	d,
	clk,
	q
	) ;

input  d;
input  clk;
inout  q;
