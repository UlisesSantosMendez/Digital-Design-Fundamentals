module comparador ( 
	a,
	b,
	x,
	y,
	z
	) ;

input [3:0] a;
input [3:0] b;
inout  x;
inout  y;
inout  z;
