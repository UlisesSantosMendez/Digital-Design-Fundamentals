module cuatrobits ( 
	clk,
	q
	) ;

input  clk;
inout [3:0] q;
