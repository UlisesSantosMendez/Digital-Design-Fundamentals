module medio ( 
	a,
	b,
	suma,
	cout
	) ;

input  a;
input  b;
inout  suma;
inout  cout;
