module mux_4 ( 
	d,
	r,
	st,
	pc,
	s,
	y
	) ;

input [3:0] d;
input [3:0] r;
input [3:0] st;
input [3:0] pc;
input [1:0] s;
inout [3:0] y;
