module display ( 
	clk,
	reset,
	d,
	q
	) ;

input  clk;
input  reset;
inout [6:0] d;
inout [3:0] q;
