module decodifdos ( 
	ra,
	rb,
	rc,
	rd,
	dispc,
	dispd,
	dispe,
	dispf
	) ;

input [3:0] ra;
input [3:0] rb;
input [3:0] rc;
input [3:0] rd;
inout [6:0] dispc;
inout [6:0] dispd;
inout [6:0] dispe;
inout [6:0] dispf;
