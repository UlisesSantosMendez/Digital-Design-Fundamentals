module decoder ( 
	a,
	d
	) ;

input [3:0] a;
inout [6:0] d;
