module c_or ( 
	a,
	d,
	c
	) ;

input  a;
input  d;
inout  c;
