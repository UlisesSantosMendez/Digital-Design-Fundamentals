module compara ( 
	a,
	b,
	z
	) ;

input [1:0] a;
input [1:0] b;
inout [1:0] z;
