module fourbits ( 
	clk,
	up,
	q
	) ;

input  clk;
input  up;
inout [3:0] q;
