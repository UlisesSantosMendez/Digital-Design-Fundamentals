module display2 ( 
	clk,
	reset,
	d
	) ;

input  clk;
input  reset;
inout [6:0] d;
