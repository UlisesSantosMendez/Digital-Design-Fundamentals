module fourbits ( 
	d,
	clk,
	clr,
	q,
	qn
	) ;

input [3:0] d;
input  clk;
input  clr;
inout [3:0] q;
inout [3:0] qn;
