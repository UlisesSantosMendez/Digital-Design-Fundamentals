module com_and ( 
	a,
	b,
	f
	) ;

input  a;
input  b;
inout  f;
