module control ( 
	clk,
	tecla,
	seg
	) ;

input  clk;
input [0:8] tecla;
inout [0:6] seg;
