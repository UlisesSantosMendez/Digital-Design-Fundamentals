module mux ( 
	a,
	b,
	c,
	d,
	s,
	z
	) ;

input [1:0] a;
input [1:0] b;
input [1:0] c;
input [1:0] d;
input [1:0] s;
inout [1:0] z;
