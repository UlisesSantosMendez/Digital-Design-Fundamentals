module mpc ( 
	cin,
	clk,
	y,
	cout,
	pc
	) ;

input  cin;
input  clk;
input [3:0] y;
inout  cout;
inout [3:0] pc;
