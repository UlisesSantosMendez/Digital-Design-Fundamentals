module comp ( 
	a,
	b,
	c
	) ;

input [1:0] a;
input [1:0] b;
inout  c;
