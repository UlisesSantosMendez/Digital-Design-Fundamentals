module contpar ( 
	p,
	clk,
	enp,
	reset,
	load,
	q
	) ;

input [3:0] p;
input  clk;
input  enp;
input  reset;
input  load;
inout [3:0] q;
