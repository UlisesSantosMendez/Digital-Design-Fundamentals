module sumador2 ( 
	cout,
	rc,
	rd,
	sum2
	) ;

inout [0:7] cout;
input [3:0] rc;
input [3:0] rd;
inout [0:7] sum2;
