module triestado ( 
	enable,
	entrada,
	salida
	) ;

input  enable;
input  entrada;
inout  salida;
