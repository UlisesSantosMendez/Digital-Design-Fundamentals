module states ( 
	clk,
	x,
	z
	) ;

input  clk;
input  x;
inout  z;
