module completo ( 
	a,
	b,
	cin,
	suma,
	cout
	) ;

input  a;
input  b;
input  cin;
inout  suma;
inout  cout;
