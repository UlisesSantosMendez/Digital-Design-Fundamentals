module ochobits ( 
	d,
	clk,
	q
	) ;

input [0:7] d;
input  clk;
inout [0:7] q;
