module sumador ( 
	a,
	b,
	suma
	) ;

input [0:3] a;
input [0:3] b;
inout [0:3] suma;
