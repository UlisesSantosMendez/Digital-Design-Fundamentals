module module ( 
	boton,
	dispa,
	dispb,
	sum
	) ;

input [0:9] boton;
inout [0:6] dispa;
inout [0:6] dispb;
inout [6:0] sum;
